CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 0 30 100 9
0 71 1536 816
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1536 816
143654930 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 784 245 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 695 388 0 1 11
0 8
0
0 0 21360 90
2 0V
11 0 25 8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 600 353 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 760 373 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 679 328 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
9 2-In AND~
219 746 287 0 3 22
0 4 5 3
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U7B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
7734 0 0
0
0
7 Pulser~
4 866 298 0 10 12
0 53 54 6 55 0 0 5 5 6
7
0
0 0 4656 512
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9914 0 0
0
0
9 2-In AND~
219 804 298 0 3 22
0 6 7 5
0
0 0 624 512
6 74LS08
-21 -24 21 -16
3 U7A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 -557942032
65 0 0 0 4 1 2 0
1 U
3747 0 0
0
0
7 Ground~
168 151 230 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
3 GND
3549 0 0
0
0
14 Logic Display~
6 888 389 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 870 388 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 852 388 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 835 389 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
10 Ascii Key~
169 524 471 0 11 12
0 25 24 23 22 56 57 58 21 0
0 53
0
0 0 4656 90
0
4 KBD3
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3363 0 0
0
0
7 74LS173
129 623 479 0 14 29
0 2 2 2 20 22 23 24 25 2
2 19 18 17 16
0
0 0 13040 692
7 74LS173
-24 -51 25 -43
2 U8
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
7 Buffer~
58 562 522 0 2 22
0 21 20
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U5C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 3 1 0
1 U
4718 0 0
0
0
7 Ground~
168 622 552 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
14 Logic Display~
6 771 156 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 753 156 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 734 156 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 717 155 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 699 155 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 682 155 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 666 155 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6843 0 0
0
0
14 Logic Display~
6 649 155 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3136 0 0
0
0
7 Ground~
168 344 343 0 1 3
0 2
0
0 0 53360 602
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
6 74LS83
105 429 352 0 14 29
0 33 32 31 30 2 2 2 2 38
34 35 36 37 59
0
0 0 13040 692
7 74LS83A
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
5670 0 0
0
0
7 Ground~
168 366 165 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6828 0 0
0
0
7 Ground~
168 266 292 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6735 0 0
0
0
7 Buffer~
58 206 252 0 2 22
0 48 47
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U5A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
8365 0 0
0
0
7 74LS193
137 787 443 0 14 29
0 10 3 11 8 19 18 17 16 60
7 15 14 13 12
0
0 0 13040 0
7 74LS193
-24 -51 25 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
4132 0 0
0
0
7 74LS273
150 575 244 0 18 37
0 9 3 34 35 36 37 39 40 41
42 33 32 31 30 29 28 27 26
0
0 0 13040 692
7 74LS273
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=20;GND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
4551 0 0
0
0
7 74LS173
129 270 226 0 14 29
0 2 2 2 47 49 50 51 52 2
2 43 44 45 46
0
0 0 13040 692
7 74LS173
-24 -51 25 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 9 10 7 11 12 13 14 1
2 6 5 4 3 15 9 10 7 11
12 13 14 1 2 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3635 0 0
0
0
6 74LS83
105 426 217 0 14 29
0 29 28 27 26 43 44 45 46 2
39 40 41 42 38
0
0 0 13040 692
7 74LS83A
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3973 0 0
0
0
10 Ascii Key~
169 160 218 0 11 12
0 52 51 50 49 61 62 63 48 0
0 54
0
0 0 4656 90
0
4 KBD1
-16 -39 12 -31
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 1 0 0 0
3 KBD
3851 0 0
0
0
74
2 0 3 0 0 12416 0 32 0 0 2 4
543 275
528 275
528 352
721 352
3 2 3 0 0 0 0 6 31 0 0 5
721 287
721 359
736 359
736 425
755 425
1 1 4 0 0 8320 0 1 6 0 0 3
785 232
766 232
766 278
3 2 5 0 0 8320 0 8 6 0 0 3
779 298
779 296
766 296
1 3 6 0 0 4224 0 8 7 0 0 2
824 289
842 289
2 10 7 0 0 8320 0 8 31 0 0 3
824 307
825 307
825 443
1 0 2 0 0 4096 0 33 0 0 65 2
238 257
238 286
4 1 8 0 0 8320 0 31 2 0 0 4
755 443
730 443
730 375
696 375
1 1 9 0 0 8320 0 32 3 0 0 3
537 284
537 340
601 340
1 1 10 0 0 8320 0 4 31 0 0 4
761 360
743 360
743 416
755 416
1 3 11 0 0 8320 0 5 31 0 0 4
680 315
666 315
666 434
749 434
14 1 12 0 0 8320 0 31 10 0 0 3
819 479
888 479
888 407
13 1 13 0 0 8320 0 31 11 0 0 3
819 470
870 470
870 406
12 1 14 0 0 8320 0 31 12 0 0 3
819 461
852 461
852 406
11 1 15 0 0 8320 0 31 13 0 0 3
819 452
835 452
835 407
14 8 16 0 0 4224 0 15 31 0 0 4
655 447
705 447
705 479
755 479
13 7 17 0 0 4224 0 15 31 0 0 4
655 456
711 456
711 470
755 470
12 6 18 0 0 4224 0 15 31 0 0 4
655 465
734 465
734 461
755 461
11 5 19 0 0 4224 0 15 31 0 0 4
655 474
726 474
726 452
755 452
1 0 2 0 0 4096 0 15 0 0 22 2
591 510
591 546
9 1 2 0 0 8192 0 15 17 0 0 3
661 510
661 546
622 546
2 1 2 0 0 4096 0 15 17 0 0 3
585 501
585 546
622 546
10 9 2 0 0 0 0 15 15 0 0 2
661 501
661 510
3 2 2 0 0 0 0 15 15 0 0 2
585 492
585 501
2 4 20 0 0 4224 0 16 15 0 0 3
577 522
577 483
591 483
8 1 21 0 0 8320 0 14 16 0 0 3
549 491
547 491
547 522
5 4 22 0 0 4224 0 15 14 0 0 4
591 474
570 474
570 467
549 467
3 6 23 0 0 4224 0 14 15 0 0 4
549 461
587 461
587 465
591 465
2 7 24 0 0 8320 0 14 15 0 0 3
549 455
549 456
591 456
1 8 25 0 0 8320 0 14 15 0 0 3
549 449
549 447
591 447
1 18 26 0 0 8320 0 18 32 0 0 3
771 174
771 203
607 203
1 0 27 0 0 8320 0 19 0 0 41 3
753 174
753 211
614 211
1 0 28 0 0 8192 0 20 0 0 40 3
734 174
734 220
619 220
1 0 29 0 0 8192 0 21 0 0 39 3
717 173
717 229
625 229
1 0 30 0 0 8192 0 22 0 0 43 3
699 173
699 239
626 239
1 0 31 0 0 4096 0 23 0 0 44 3
682 173
682 248
619 248
1 0 32 0 0 4096 0 24 0 0 45 3
666 173
666 259
614 259
1 0 33 0 0 4096 0 25 0 0 46 3
649 173
649 273
607 273
1 15 29 0 0 20608 0 34 32 0 0 8
394 257
382 257
382 278
483 278
483 174
625 174
625 230
607 230
2 16 28 0 0 20608 0 34 32 0 0 8
394 248
371 248
371 291
487 291
487 179
619 179
619 221
607 221
3 17 27 0 0 0 0 34 32 0 0 8
394 239
365 239
365 295
491 295
491 183
614 183
614 212
607 212
4 18 26 0 0 0 0 34 32 0 0 7
394 230
360 230
360 299
497 299
497 188
607 188
607 203
4 14 30 0 0 12416 0 27 32 0 0 8
397 365
373 365
373 430
575 430
575 324
626 324
626 239
607 239
3 13 31 0 0 12416 0 27 32 0 0 8
397 374
379 374
379 424
569 424
569 318
619 318
619 248
607 248
2 12 32 0 0 12416 0 27 32 0 0 8
397 383
385 383
385 419
563 419
563 314
614 314
614 257
607 257
1 11 33 0 0 12416 0 27 32 0 0 7
397 392
391 392
391 413
556 413
556 309
607 309
607 266
10 3 34 0 0 8320 0 27 32 0 0 4
461 365
522 365
522 266
543 266
11 4 35 0 0 8320 0 27 32 0 0 4
461 356
515 356
515 257
543 257
12 5 36 0 0 8320 0 27 32 0 0 4
461 347
508 347
508 248
543 248
13 6 37 0 0 8320 0 27 32 0 0 4
461 338
502 338
502 239
543 239
6 0 2 0 0 4224 0 27 0 0 52 2
397 347
351 347
5 1 2 0 0 0 0 27 26 0 0 3
397 356
351 356
351 344
7 0 2 0 0 0 0 27 0 0 54 2
397 338
351 338
8 1 2 0 0 0 0 27 26 0 0 3
397 329
351 329
351 344
14 9 38 0 0 8320 0 34 27 0 0 5
458 176
478 176
478 283
397 283
397 311
10 7 39 0 0 4224 0 34 32 0 0 2
458 230
543 230
11 8 40 0 0 4224 0 34 32 0 0 2
458 221
543 221
12 9 41 0 0 4224 0 34 32 0 0 2
458 212
543 212
13 10 42 0 0 4224 0 34 32 0 0 2
458 203
543 203
1 9 2 0 0 0 0 28 34 0 0 3
366 159
394 159
394 176
11 5 43 0 0 4224 0 33 34 0 0 2
302 221
394 221
12 6 44 0 0 4224 0 33 34 0 0 2
302 212
394 212
13 7 45 0 0 4224 0 33 34 0 0 2
302 203
394 203
14 8 46 0 0 4224 0 33 34 0 0 2
302 194
394 194
2 1 2 0 0 0 0 33 29 0 0 3
232 248
232 286
266 286
9 1 2 0 0 0 0 33 29 0 0 3
308 257
308 286
266 286
10 9 2 0 0 0 0 33 33 0 0 2
308 248
308 257
3 2 2 0 0 0 0 33 33 0 0 2
232 239
232 248
4 2 47 0 0 8320 0 33 30 0 0 3
238 230
221 230
221 252
8 1 48 0 0 8320 0 35 30 0 0 3
185 238
191 238
191 252
4 5 49 0 0 4224 0 35 33 0 0 4
185 214
222 214
222 221
238 221
3 6 50 0 0 4224 0 35 33 0 0 4
185 208
227 208
227 212
238 212
2 7 51 0 0 8320 0 35 33 0 0 3
185 202
185 203
238 203
1 8 52 0 0 8320 0 35 33 0 0 3
185 196
185 194
238 194
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
